
`timescale 1 ns/10 ps  // time-unit = 1 ns, precision = 10 ps

module bf16_unit_tb();

	localparam period = 10; // 10 ns


	integer i;
	integer j;
	integer k;
	
	reg clk; 
	reg reset;
	reg [15:0] in1; 
	reg [15:0] in2;
	reg [15:0] in3;
	reg [15:0] in4; 
	reg [15:0] in5;
	reg [15:0] in6;
	reg [15:0] in7; 
	reg [15:0] in8;
	reg [15:0] in9;
	reg [15:0] in10; 
	reg [15:0] in11;
	reg [15:0] in12;
	reg [15:0] in13; 
	reg [15:0] in14;
	reg [15:0] in15;
	reg [15:0] in16;
	reg [15:0] in17;
	reg [15:0] in18; 
	reg [4:0] funct5;
	wire [15:0] result;
	
	bf16_unit UUT(.clk(clk), 
				  .reset(reset), 
				  .in1(in1),
				  .in2(in2),
				  .in3(in3),
				  .in4(in4),
				  .in5(in5),
				  .in6(in6),
				  .in7(in7),
				  .in8(in8),
				  .in9(in9),
				  .in10(in10),
				  .in11(in11),
				  .in12(in12),
				  .in13(in13),
				  .in14(in14),
				  .in15(in15),
				  .in16(in16),
				  .in17(in17),
				  .in18(in18),
				  .funct5(funct5),
				  .result(result) );
				  

	  // generate the clock
	  initial begin
		clk = 1'b1;
		forever #5 clk = ~clk;
	  end
	  
	  // Generate the reset
	  initial begin
	   reset = 1'b0;
	   #15
	   reset = 1'b1;
	  end
	  
	  // Generate funct5
	  initial begin
	  	  funct5 = 0; 
	  	  #40
	      #200 funct5 = 5'b00001; 
	      #200 funct5 = 5'b00010; 
	      #200 funct5 = 5'b00100; 
	      #200 funct5 = 5'b00101;
	      #200 funct5 = 5'b00111;  
	  end
	  
	  // Generate in1
	  initial begin
	  	  in1 = 16'b0000000000000000;
	  	  #30
	      for (i = 0; i < 6; i = i+1) begin
	  		  #10 in1 = 16'b0100010001011000;
	          #10 in1 = 16'b1100010001111000;
              #10 in1 = 16'b0001010001000010;
              #10 in1 = 16'b0100101001001011;
              #10 in1 = 16'b1000000011101000;
              #10 in1 = 16'b0111111110011000;
	          #10 in1 = 16'b1100011001001101;
	          #10 in1 = 16'b1000000001001101;
	          #10 in1 = 16'b0000000000000000; 
	          #10 in1 = 16'b1111111110000000; 
              #10 in1 = 16'b0100000011110011; 
              #10 in1 = 16'b1100000011110011; 
              #10 in1 = 16'b0100001100101100; 
              #10 in1 = 16'b0100001100001100; 
              #10 in1 = 16'b0100001101101100; 
              #10 in1 = 16'b1011111010000000; 
              #10 in1 = 16'b1100000011000000; 
              #10 in1 = 16'b0010101010000111; 
              #10 in1 = 16'b0010101010000111; 
              #10 in1 = 16'b0100010110100000;
          end
      end
	  
	  // Generate in2
	  initial begin
	  	  in2 = 16'b0000000000000000;
	  	  #30
	      for (j = 0; j < 6; j = j+1) begin
	  		  #10 in2 = 16'b1100010001111000;
	          #10 in2 = 16'b0100010001011000;
              #10 in2 = 16'b0001011001001011;
              #10 in2 = 16'b0000001001101000;
              #10 in2 = 16'b0000001001101000;
              #10 in2 = 16'b1000100101001000;
	          #10 in2 = 16'b1100011110011000;
	          #10 in2 = 16'b1000000100001010;
	          #10 in2 = 16'b0000000000011100; 
	          #10 in2 = 16'b0100000011110011; 
              #10 in2 = 16'b0100000011110011; 
              #10 in2 = 16'b0100000011110011; 
              #10 in2 = 16'b1100010111101010; 
              #10 in2 = 16'b1100001101101010; 
              #10 in2 = 16'b1100001101101010; 
              #10 in2 = 16'b0100000011000000; 
              #10 in2 = 16'b1100000111001000; 
              #10 in2 = 16'b0110101010100111; 
              #10 in2 = 16'b0100010000100011; 
              #10 in2 = 16'b0100000110100000;
          end
      end
      
      // Generate in3
	  initial begin
	  	  in3 = 16'b0000000000000000;
	  	  #30
	      for (k = 0; k < 6; k = k+1) begin
	  		  #10 in3 = 16'b1100010001111000;
	          #10 in3 = 16'b0100010001011000;
              #10 in3 = 16'b0001011001001011;
              #10 in3 = 16'b0000001001101000;
              #10 in3 = 16'b0000001001101000;
              #10 in3 = 16'b1000100101001000;
	          #10 in3 = 16'b1100011110011000;
	          #10 in3 = 16'b1000000100001010;
	          #10 in3 = 16'b0000000000011100; 
	          #10 in3 = 16'b0100000011110011; 
              #10 in3 = 16'b0100000011110011; 
              #10 in3 = 16'b0100000011110011; 
              #10 in3 = 16'b1100010111101010; 
              #10 in3 = 16'b1100001101101010; 
              #10 in3 = 16'b1100001101101010; 
              #10 in3 = 16'b0100000011000000; 
              #10 in3 = 16'b1100000111001000; 
              #10 in3 = 16'b0110101010100111; 
              #10 in3 = 16'b0100010000100011; 
              #10 in3 = 16'b0100000110100000;
          end
      end
	  
	  // Generate in1
	  initial begin
	  	  #1500
	  	  in1 = 16'b0011110111111000;
	  	  #10
	  	  in1 = 16'b0100000001100000;
	  end
	  
	  // Generate in2
	  initial begin
	  	  #1500
	  	  in2 = 16'b0011110101010101;
	  	  #10
	  	  in2 = 16'b0100000100010000;
	  end
	  
	  // Generate in3
	  initial begin
	  	  #1500
	  	  in3 = 16'b0011110111111100;
	  	  #10
	  	  in3 = 16'b0100000000110000;
	  end
	  
	  // Generate in4
	  initial begin
	  	  in4 = 16'b0000000000000000;
	  	  #1500
	  	  in4 = 16'b0011111101011010;
	  	  #10
	  	  in4 = 16'b0011111110000000;
	  end
	  
	  // Generate in5
	  initial begin
	  	  in5 = 16'b0000000000000000;
	  	  #1500
	  	  in5 = 16'b0011111100011001;
	  	  #10
	  	  in5 = 16'b0011111110000000;
	  end
	  
	  // Generate in6
	  initial begin
	  	  in6 = 16'b0000000000000000;
	  	  #1500
	  	  in6 = 16'b0011111010101000;
	  	  #10
	  	  in6 = 16'b0011111110000000;
	  end
	  
	  // Generate in7
	  initial begin
	  	  in7 = 16'b0000000000000000;
	  	  #1500
	  	  in7 = 16'b0000000000000000;
	  	  #10
	  	  in7 = 16'b0011111110000000;
	  end
	  
	  // Generate in8
	  initial begin
	  	  in8 = 16'b0000000000000000;
	  	  #1500
	  	  in8 = 16'b0000000000000000;
	  	  #10
	  	  in8 = 16'b0011111110000000;
	  end
	  
	  // Generate in9
	  initial begin
	  	  in9 = 16'b0000000000000000;
	  	  #1500
	  	  in9 = 16'b0000000000000000;
	  	  #10
	  	  in9 = 16'b0011111110000000;
	  end
	  
	  // Generate in10
	  initial begin
	  	  in10 = 16'b0000000000000000;
	  	  #1500
	  	  in10 = 16'b0000000000000000;
	  	  #10
	  	  in10 = 16'b0011111110000000;
	  end
	  
	  // Generate in11
	  initial begin
	  	  in11 = 16'b0000000000000000;
	  	  #1500
	  	  in11 = 16'b0000000000000000;
	  	  #10
	  	  in11 = 16'b0011111110000000;
	  end
	  
	  // Generate in12
	  initial begin
	  	  in12 = 16'b0000000000000000;
	  	  #1500
	  	  in12 = 16'b0000000000000000;
	  	  #10
	  	  in12 = 16'b0011111110000000;
	  end
	  
	  // Generate in13
	  initial begin
	  	  in13 = 16'b0000000000000000;
	  	  #1500
	  	  in13 = 16'b0000000000000000;
	  	  #10
	  	  in13 = 16'b0011111110000000;
	  end
	  
	  // Generate in14
	  initial begin
	  	  in14 = 16'b0000000000000000;
	  	  #1500
	  	  in14 = 16'b0000000000000000;
	  	  #10
	  	  in14 = 16'b0011111110000000;
	  	  #10
	  	  in14 = 16'b0100000000000000;
	  end
	  
	  // Generate in15
	  initial begin
	  	  in15 = 16'b0000000000000000;
	  	  #1500
	  	  in15 = 16'b0000000000000000;
	  	  #10
	  	  in15 = 16'b0011111110000000;
	  end
	  
	  // Generate in16
	  initial begin
	  	  in16 = 16'b0000000000000000;
	  	  #1500
	  	  in16 = 16'b0000000000000000;
	  	  #10
	  	  in16 = 16'b0011111110000000;
	  	  #10
	  	  in16 = 16'b0100000000000000;
	  end
	  
	  // Generate in17
	  initial begin
	  	  in17 = 16'b0000000000000000;
	  	  #1500
	  	  in17 = 16'b0000000000000000;
	  	  #10
	  	  in17 = 16'b0011111110000000;
	  	  #10
	  	  in17 = 16'b0100000000000000;
	  end
	  
	  // Generate in18
	  initial begin
	  	  in18 = 16'b0000000000000000;
	  	  #1500
	  	  in18 = 16'b0000000000000000;
	  	  #10
	  	  in18 = 16'b0011111110000000;
	  	  #10
	  	  in18 = 16'b0100000000000000;
	  end

endmodule
