
`timescale 1 ns/10 ps  // time-unit = 1 ns, precision = 10 ps

module bf16_unit_tb();

	localparam period = 10; // 10 ns

	integer i;
	integer m;
	integer k;
	integer l;

	reg clk; 
	reg reset;
	reg [15:0] in1; 
	reg [15:0] in2;
	reg [15:0] in3; 
	reg [4:0] funct5;
	wire [15:0] result;
	
	bf16_unitt UUT(.clk(clk), 
		.reset(reset), 
		.in1(in1),
		.in2(in2),
		.in3(in3),
		.funct5(funct5),
		.result(result) );
				  

	// generate the clock
	initial begin
		clk = 1'b1;
		forever #5 clk = ~clk;
	end
	
	// Generate the reset
	initial begin
		reset = 1'b0;
		#15
		reset = 1'b1;
	end
	
	// Generate funct5
	initial begin
		funct5 = 0; 
		#40
		for (i = 0; i < 2; i = i+1) begin
			#200 funct5 = i + 1; 
		end
	end
	
	// Generate in1
	initial begin
		in1 = 16'b0000000000000000;
		#30
		for (k = 0; k < 3; k = k+1) begin
			#10 in1 = 16'b0100010001011000; 
			#10 in1 = 16'b1100010001111000; 
			#10 in1 = 16'b0001010001000010;
			#10 in1 = 16'b0100101001001011; 
			#10 in1 = 16'b1000000011101000; 
			#10 in1 = 16'b0111111110011000; 
			#10 in1 = 16'b1100011001001101; 
			#10 in1 = 16'b1000000001001101; 
			#10 in1 = 16'b0000000000000000; 
			#10 in1 = 16'b1111111110000000; 
			#10 in1 = 16'b0100000011110011; 
			#10 in1 = 16'b1100000011110011; 
			#10 in1 = 16'b0100001100101100; 
			#10 in1 = 16'b0100001100001100; 
			#10 in1 = 16'b0100001101101100; 
			#10 in1 = 16'b1011111010000000; 
			#10 in1 = 16'b1100000011000000; 
			#10 in1 = 16'b0010101010000111; 
			#10 in1 = 16'b0010101010000111; 
			#10 in1 = 16'b0100010110100000; 
		end
	end
	
	// Generate in2
	initial begin
		in2 = 16'b0000000000000000;
		#30
		for (m = 0; m < 3; m = m+1) begin
			#10 in2 = 16'b1100010001111000;
			#10 in2 = 16'b0100010001011000;
			#10 in2 = 16'b0001011001001011;
			#10 in2 = 16'b0000001001101000;
			#10 in2 = 16'b0000001001101000;
			#10 in2 = 16'b1000100101001000;
			#10 in2 = 16'b1100011110011000;
			#10 in2 = 16'b1000000100001010;
			#10 in2 = 16'b0000000000011100; 
			#10 in2 = 16'b0100000011110011; 
			#10 in2 = 16'b0100000011110011; 
			#10 in2 = 16'b0100000011110011; 
			#10 in2 = 16'b1100010111101010; 
			#10 in2 = 16'b1100001101101010; 
			#10 in2 = 16'b1100001101101010; 
			#10 in2 = 16'b0100000011000000; 
			#10 in2 = 16'b1100000111001000; 
			#10 in2 = 16'b0110101010100111; 
			#10 in2 = 16'b0100010000100011; 
			#10 in2 = 16'b0100000110100000;
		end
	end
      
	// Generate in3
	initial begin
		in3 = 16'b0000000000000000;
		#30
		for (l = 0; l < 3; l = l+1) begin
			#10 in3 = 16'b1100010001111000;
			#10 in3 = 16'b0100010001011000;
			#10 in3 = 16'b0001011001001011;
			#10 in3 = 16'b0000001001101000;
			#10 in3 = 16'b0000001001101000;
			#10 in3 = 16'b1000100101001000;
			#10 in3 = 16'b1100011110011000;
			#10 in3 = 16'b1000000100001010;
			#10 in3 = 16'b0000000000011100; 
			#10 in3 = 16'b0100000011110011; 
			#10 in3 = 16'b0100000011110011; 
			#10 in3 = 16'b0100000011110011; 
			#10 in3 = 16'b1100010111101010; 
			#10 in3 = 16'b1100001101101010; 
			#10 in3 = 16'b1100001101101010; 
			#10 in3 = 16'b0100000011000000; 
			#10 in3 = 16'b1100000111001000; 
			#10 in3 = 16'b0110101010100111; 
			#10 in3 = 16'b0100010000100011; 
			#10 in3 = 16'b0100000110100000;
		end
	end

endmodule
